-------------------------------------------------------------------------------
--                                                                      
--                        Counter Project Base
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         io_ctrl
--
-- FILENAME:       io_ctrl_rtl.vhd
-- 
-- ARCHITECTURE:   RTL
-- 
-- ENGINEER:       <>
--
-- DATE:           <>
--
-- VERSION:        <>
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This describes the architecture of the io control sub unit
--                 of the counter VHDL class example.
--
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------
--                                                                      
-- CHANGES:
--                 1.0 - initial version
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
-- do NOT use std_logic_arith
library work;
use work.counter_util_pkg.all;
use work.counter_comp_pkg.all;

architecture rtl of io_ctrl is

begin

end rtl;
